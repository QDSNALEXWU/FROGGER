module digitfont( input logic Clk,
               	// from right to left
               	input logic [0:3] digit,  	
						output logic [0:13][0:13][0:5] font 
				  );


logic [0:13][0:13][0:5] zero_font ;  
logic [0:13][0:13][0:5] one_font ; 
logic [0:13][0:13][0:5] two_font ; 
logic [0:13][0:13][0:5] three_font ;  
logic [0:13][0:13][0:5] four_font ;  
logic [0:13][0:13][0:5] five_font ; 
logic [0:13][0:13][0:5] six_font ;
logic [0:13][0:13][0:5] seven_font ; 
logic [0:13][0:13][0:5] eight_font ; 
logic [0:13][0:13][0:5] nine_font ; 



// assign the font values
always_comb
begin
	zero_font <= '{
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{0, 0, 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	'{0, 0, 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	'{0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }
	};

	one_font<='{
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }
	};

	two_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }
	};

	three_font<='{
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	four_font<='{
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }
	};


	five_font<='{
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};


	six_font<='{
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	seven_font<='{
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }
	};

	eight_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2 },  
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2 },   
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }, 
	'{ 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	nine_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }
	};
end 

//output the value

always_comb
begin
	case (digit)
		4'b0000 : 
			begin 	
				font = zero_font ; 
			end	
		
		4'b0001 : 
			begin 	
				font = one_font ; 
			end	

		4'b0010 : 
			begin 	
				font = two_font ; 
			end	

		4'b0011  : 
			begin 	
				font = three_font ; 
			end		

		4'b0100 : 
			begin 	
				font = four_font ; 
			end		

		4'b0101 : 
			begin 	
				font = five_font ; 
			end	

		4'b0110 : 
			begin 	
				font = six_font ; 
			end

		4'b0111 : 
			begin 	
				font = seven_font ; 
			end		

		4'b1000: 
			begin 	
				font = eight_font ; 
			end	
		
		4'b1001 : 
			begin 	
				font = nine_font ; 
			end	

		default : 
			begin      
				font = zero_font ; 
			end 	
		
	endcase	



end

endmodule


