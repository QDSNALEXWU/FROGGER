module lab8( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK      //SDRAM Clock
                    );
    
    // ********* self-delcrared varibales **********************
    // ********* VARIABLES GROUP 1 ***************************** 
    logic [0:5] colorcode;
    logic [0:15][0:16][0:5] frog_font ;
    logic [0:15][0:24][0:5] firetruck_font ;
    logic [0:13][0:18][0:5] bus_font ;
    logic [0:15][0:22][0:5] motorcycle_font ;
    logic [0:15][0:26][0:5] shortlog_font ;
    logic [0:15][0:49][0:5] mediumlog_font ;
    logic [0:15][0:72][0:5] longlog_font ; 
    logic [0:11][0:13][0:5] heart_font ;
    logic [0:15][0:15][0:5] Oneshell_font ;
    logic [0:15][0:32][0:5] Twoshell_font ;
    logic [0:15][0:49][0:5] Threeshell_font ; 
    logic [0:12][0:26][0:5] gator_font ;
    logic [0:23][0:26][0:5] vader_font ; 
    logic [0:11][0:27][0:5] policecar_font ;
	logic [0:13][0:24][0:5] truck_font ;   	
    logic [0:17][0:22][0:5] skull_font ;
    logic [0:13][0:13][0:5] S_font ;  
    logic [0:13][0:13][0:5] C_font ;  
    logic [0:13][0:13][0:5] O_font ; 
    logic [0:13][0:13][0:5] R_font ;  
    logic [0:13][0:13][0:5] E_font ;  
    logic [0:13][0:13][0:5] T_font ;  
    logic [0:13][0:13][0:5] I_font ;
    logic [0:13][0:13][0:5] M_font ; 
    logic [3:0]  ten ;  
    logic [3:0]  hundred ;
    logic [3:0]  thousand ; 

    
	 // ********* VARIABLES GROUP 2 *****************************     
    logic Reset_h, Clk;
    logic [15:0] keycode;
    
    assign Clk = CLOCK_50;
    assign {Reset_h} = ~(KEY[0]);  // The push buttons are active low
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w,hpi_cs;
    


    // Self Declared Variables
    logic [9:0] DrawX,DrawY,BallX,BallY,BallS;

    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),    
                            .OTG_RST_N(OTG_RST_N)
    );
     
     //The connections for nios_system might be named different depending on how you set up Qsys
     nios_system nios_system_unit(
                             .clk_clk(Clk),         
                             .reset_reset_n(KEY[0]),   
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w)
    );
    
     //Fill in the connections for the rest of the modules 
    
	 // interaction with VGA 
     VGA_controller vga_controller_instance( .* , .Reset(Reset_h) );
    
	 // keyboard input handler  
	 ball ball_instance( .*, .Reset(~KEY[2]), .frame_clk(VGA_VS));  
    
	 // store all the font we need 
	 fontawesome fontawesome_instance(.*);
    
     // get all the text_font
     letterfont letterfont_instance(.*);

	 // game logic control unit 
	 frogger_game game_instance(.*);
    
	 // map RGB value with color code 
	 color_mapper color_instance(.*);
    
     HexDriver hex_inst_0 (keycode[3:0], HEX0);
     HexDriver hex_inst_1 (keycode[7:4], HEX1);

endmodule
