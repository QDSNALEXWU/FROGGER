module fontawesome(input logic Clk,
                   // Y X L 
                   output logic [0:15][0:16][0:5] frog_font,
                   output logic [0:15][0:24][0:5] firetruck_font,
                   output logic [0:13][0:18][0:5] bus_font,
                   output logic [0:15][0:22][0:5] motorcycle_font,
                   output logic [0:8][0:26][0:5] shortlog_font,
                   output logic [0:8][0:49][0:5] mediumlog_font,
                   output logic [0:8][0:72][0:5] longlog_font,
                   output logic [0:15][0:7][0:5] heart_font 
                  );

						
always_comb
    begin
  
      // frog font 17 x 16 
      frog_font <= '{ 
      '{ 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0 }, 
      '{ 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0 },  
      '{ 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0 },
      '{ 0, 1, 0, 1, 1, 0, 0, 2, 2, 2, 0, 0, 1, 1, 0, 1, 0 },
      '{ 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0 },
      '{ 0, 0, 1, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 0, 1, 0, 0 },
      '{ 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0 },
      '{ 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 2, 1 },
      '{ 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 1 },
      '{ 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0 },
      '{ 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0 },
      '{ 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0 },
      '{ 0, 1, 1, 2, 2, 2, 2, 2, 0, 2, 2, 2, 2, 2, 1, 1, 0 },
      '{ 1, 2, 1, 2, 2, 2, 2, 0, 0, 0, 2, 2, 2, 2, 1, 2, 1 },
      '{ 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1 },
      '{ 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0 }
      } ;

      // fire truck font 25 x 16
      firetruck_font <=  '{ 
      '{ 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
      '{ 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
      '{ 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 }, 
      '{ 0, 0, 3, 4, 4, 4, 3, 3, 4, 4, 3, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1 }, 
      '{ 0, 3, 3, 4, 4, 4, 3, 3, 4, 4, 3, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 },
      '{ 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0 },
      '{ 0, 3, 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0 },
      '{ 0, 3, 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 6, 6, 6, 3, 6, 6, 6, 3, 6, 6, 6, 3, 0 }, 
      '{ 0, 3, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 6, 6, 6, 3, 6, 3, 3, 3, 3, 3, 6, 3, 3 }, 
      '{ 0, 3, 6, 6, 3, 1, 1, 1, 1, 3, 3, 3, 6, 6, 6, 3, 3, 1, 1, 1, 1, 3, 3, 3, 3 },
      '{ 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 7, 7, 7 }, 
      '{ 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7 },
      '{ 0, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7 }, 
      '{ 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 ,0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0 ,0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0 }
      };

      // Bus font 19 x 14
      bus_font <= '{
      '{ 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0 },
      '{ 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 3, 3, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3 },
      '{ 3, 3, 3, 6, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3 },
      '{ 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 }, 
      '{ 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 6, 3, 6, 6, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 3 },
      '{ 6, 3, 6, 6, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 3 },
      '{ 3, 3, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 5, 3, 3, 3, 3, 1, 1, 3, 3, 3, 3, 3, 3, 1, 1, 3, 3, 5, 3 },
      '{ 3, 3, 3, 3, 1, 4, 4, 1, 3, 3, 3, 3, 1, 4, 4, 1, 3, 3, 3 }, 
      '{ 0, 0, 0, 0, 1, 4, 4, 0, 0, 0, 0, 0, 1, 4, 4, 1, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0 }
      };

      // Motorcycle font 23 x 16
      motorcycle_font <= '{
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 5, 5, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 5, 5, 5, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 5, 5, 5, 5, 5, 1, 1, 1, 1, 1, 1, 1, 1, 0 },
      '{ 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 3, 3, 3, 3, 3, 3, 3, 1 },
      '{ 0, 1, 1, 1, 1, 1, 1, 1, 1, 6, 6, 6, 6, 6, 6, 1, 1, 1, 1, 1, 1, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 0, 1, 6, 6, 6, 6, 6, 1, 0, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 6, 6, 6, 6, 1, 1, 0, 0, 0, 0, 0, 1, 0 },
      '{ 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 6, 6, 6, 1, 1, 1, 0, 1, 0, 0, 0, 1 }, 
      '{ 1, 0, 0, 1, 5, 1, 0, 0, 1, 0, 1, 6, 6, 6, 1, 0, 0, 1, 5, 1, 0, 0, 1 }, 
      '{ 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1 },
      '{ 1, 0, 0, 1, 5, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 5, 1, 0, 0, 1 },
      '{ 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1 },
      '{ 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0 }
      };


       // Short Log (27 x 9)
      shortlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };

       // Medium Log (50 x 9)
       mediumlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };


       // Long Log (73 x 9) 
       longlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };

      // Heart  8x16 
      heart_font <= '{
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 0
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 1
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 2
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 3
        '{ 0, 1, 1, 0, 1, 1, 0, 0 }, // 4  ** **
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 5 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 6 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 7 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 8 *******
        '{ 0, 1, 1, 1, 1, 1, 0, 0 }, // 9  *****
        '{ 0, 0, 1, 1, 1, 0, 0, 0 }, // a   ***
        '{ 0, 0, 0, 1, 0, 0, 0, 0 }, // b    *
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // c
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // d
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // e
        '{ 0, 0, 0, 0, 0, 0, 0, 0 } // f
    };
	end
endmodule

