module fontawesome(input logic Clk,
                   // Y X L 
                   output logic [0:15][0:16][0:5] frog_font,
                   output logic [0:15][0:24][0:5] firetruck_font,
                   output logic [0:13][0:18][0:5] bus_font,
                   output logic [0:15][0:22][0:5] motorcycle_font,
                   output logic [0:8][0:26][0:5] shortlog_font,
                   output logic [0:8][0:49][0:5] mediumlog_font,
                   output logic [0:8][0:72][0:5] longlog_font,
                   output logic [0:15][0:7][0:5] heart_font, 
						 output logic [0:15][0:15][0:5] Oneshell_font,
						 output logic [0:15][0:32][0:5] Twoshell_font,
						 output logic [0:15][0:49][0:5] Threeshell_font,  
                   output logic [0:12][0:26][0:5] gator_font,
                   output logic [0:23][0:26][0:5] vader_font, 
						 output logic [0:11][0:27][0:5] policecar_font,
						 output logic [0:13][0:24][0:5] truck_font,   	
					    output logic [0:17][0:22][0:5] skull_font	
						);
						
always_comb
    begin
  
      // frog font 17 x 16 
      frog_font <= '{ 
      '{ 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0 }, 
      '{ 0, 0, 1, 11, 11, 11, 1, 0, 0, 0, 1, 11, 11, 11, 1, 0, 0 },  
      '{ 0, 1, 11, 1, 1, 11, 11, 1, 1, 1, 11, 11, 1, 1, 11, 1, 0 },
      '{ 0, 1, 11, 1, 1, 11, 11, 2, 2, 2, 11, 11, 1, 1, 11, 1, 0 },
      '{ 0, 1, 11, 11, 11, 11, 11, 2, 2, 2, 11, 11, 11, 11, 11, 1, 0 },
      '{ 0, 0, 1, 11, 11, 11, 2, 2, 2, 2, 2, 11, 11, 11, 1, 0, 0 },
      '{ 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0 },
      '{ 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 2, 1 },
      '{ 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 1 },
      '{ 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0 },
      '{ 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0 },
      '{ 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0 },
      '{ 0, 1, 1, 2, 2, 2, 2, 2, 11, 2, 2, 2, 2, 2, 1, 1, 0 },
      '{ 1, 2, 1, 2, 2, 2, 2, 11, 11, 11, 2, 2, 2, 2, 1, 2, 1 },
      '{ 1, 2, 2, 2, 1, 2, 1, 11, 11, 11, 1, 2, 1, 2, 2, 2, 1 },
      '{ 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0 }
      } ;

      // fire truck font 25 x 16
      firetruck_font <=  '{ 
      '{ 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
      '{ 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
      '{ 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 }, 
      '{ 0, 0, 3, 4, 4, 4, 3, 3, 4, 4, 3, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1 }, 
      '{ 0, 3, 3, 4, 4, 4, 3, 3, 4, 4, 3, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 },
      '{ 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0 },
      '{ 0, 3, 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0 },
      '{ 0, 3, 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 6, 6, 6, 3, 6, 6, 6, 3, 6, 6, 6, 3, 0 }, 
      '{ 0, 3, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 6, 6, 6, 3, 6, 3, 3, 3, 3, 3, 6, 3, 3 }, 
      '{ 0, 3, 6, 6, 3, 1, 1, 1, 1, 3, 3, 3, 6, 6, 6, 3, 3, 1, 1, 1, 1, 3, 3, 3, 3 },
      '{ 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 7, 7, 7 }, 
      '{ 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7 },
      '{ 0, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7, 7, 7, 7, 1, 1, 6, 6, 1, 1, 7, 7, 7 }, 
      '{ 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 ,0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0 ,0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0 }
      };

      // Bus font 19 x 14
      bus_font <= '{
      '{ 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0 },
      '{ 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 3, 3, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3 },
      '{ 3, 3, 3, 6, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3 },
      '{ 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 }, 
      '{ 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 6, 3, 6, 6, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 3 },
      '{ 6, 3, 6, 6, 3, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 6, 6, 3, 3 },
      '{ 3, 3, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 },
      '{ 5, 3, 3, 3, 3, 1, 1, 3, 3, 3, 3, 3, 3, 1, 1, 3, 3, 5, 3 },
      '{ 3, 3, 3, 3, 1, 4, 4, 1, 3, 3, 3, 3, 1, 4, 4, 1, 3, 3, 3 }, 
      '{ 0, 0, 0, 0, 1, 4, 4, 0, 0, 0, 0, 0, 1, 4, 4, 1, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0 }
      };

      // Motorcycle font 23 x 16
      motorcycle_font <= '{
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 5, 5, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 5, 5, 5, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 5, 5, 5, 5, 5, 1, 1, 1, 1, 1, 1, 1, 1, 0 },
      '{ 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 3, 3, 3, 3, 3, 3, 3, 1 },
      '{ 0, 1, 1, 1, 1, 1, 1, 1, 1, 6, 6, 6, 6, 6, 6, 1, 1, 1, 1, 1, 1, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 0, 1, 6, 6, 6, 6, 6, 1, 0, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 6, 6, 6, 6, 1, 1, 0, 0, 0, 0, 0, 1, 0 },
      '{ 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 6, 6, 6, 1, 1, 1, 0, 1, 0, 0, 0, 1 }, 
      '{ 1, 0, 0, 1, 5, 1, 0, 0, 1, 0, 1, 6, 6, 6, 1, 0, 0, 1, 5, 1, 0, 0, 1 }, 
      '{ 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1 },
      '{ 1, 0, 0, 1, 5, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 5, 1, 0, 0, 1 },
      '{ 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1 },
      '{ 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0 }
      };


       // Short Log (27 x 9)
      shortlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };

       // Medium Log (50 x 9)
       mediumlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };


       // Long Log (73 x 9) 
       longlog_font <= '{
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 1, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 1, 1, 0, 1 }, 
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 8, 8, 8, 1, 1, 1, 8, 8, 8, 8, 8, 8, 8, 1, 1, 8, 8, 8, 8, 8, 1, 0, 0, 0, 0, 1 },
      '{ 0, 1, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0, 0, 1, 0 },
      '{ 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }
      };

      // Heart  8x16 
      heart_font <= '{
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 0
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 1
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 2
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // 3
        '{ 0, 1, 1, 0, 1, 1, 0, 0 }, // 4  ** **
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 5 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 6 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 7 *******
        '{ 1, 1, 1, 1, 1, 1, 1, 0 }, // 8 *******
        '{ 0, 1, 1, 1, 1, 1, 0, 0 }, // 9  *****
        '{ 0, 0, 1, 1, 1, 0, 0, 0 }, // a   ***
        '{ 0, 0, 0, 1, 0, 0, 0, 0 }, // b    *
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // c
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // d
        '{ 0, 0, 0, 0, 0, 0, 0, 0 }, // e
        '{ 0, 0, 0, 0, 0, 0, 0, 0 } // f
    };


     // gator 27x13 
     gator_font <= '{
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2 }, 
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 2, 12, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 2 },
      '{ 0, 0, 0, 0, 0, 0, 2, 12, 1, 1, 12, 1, 0, 0, 2, 0, 2, 0, 2, 0, 0, 0, 0, 0, 2, 12, 2 }, 
      '{ 0, 0, 0, 0, 0, 0, 2, 12, 11, 1, 12, 12, 2, 2, 12, 2, 12, 2, 12, 2, 0, 0, 0, 2, 12, 12, 2 }, 
      '{ 0, 2, 2, 2, 0, 2, 12, 12, 12, 12, 12, 12, 2, 12, 12, 12, 12, 12, 12, 12, 2, 2, 2, 12, 12, 2, 0 }, 
      '{ 2, 12, 1, 12, 2, 12, 12, 12, 12, 12, 12, 12, 12, 12, 2, 2, 12, 2, 2, 12, 12, 12, 12, 12, 12, 2, 0 },
      '{ 2, 12, 12, 12, 12, 12, 12, 2, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 2, 0, 0 },
      '{ 0, 2, 2, 2, 2, 2, 2, 12, 12, 12, 12, 12, 2, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 2, 0, 0, 0 }, 
      '{ 0, 0, 2, 12, 12, 12, 12, 12, 12, 12, 12, 2, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 1, 0, 0, 0, 0 }, 
      '{ 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 2, 2, 2, 0, 2, 2, 2, 2, 12, 12, 2, 0, 0, 0 }, 
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 2, 0, 2, 12, 2, 2, 12, 2, 12, 12, 1, 0, 0, 0 }, 
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 2, 2, 2, 2, 0, 2, 2, 0, 0, 0, 0 }
     };


    // vader 27x24
     vader_font <= '{
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 6, 1, 6, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 1, 1, 1, 1, 6, 6, 6, 6, 6, 1, 6, 6, 6, 6, 6, 1, 1, 1, 1, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 1, 1, 1, 6, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 6, 1, 1, 1, 0, 0, 0, 0 },
      '{ 0, 0, 0, 0, 1, 1, 6, 6, 1, 1, 1, 1, 1, 6, 1, 1, 1, 1, 1, 6, 6, 1, 1, 0, 0, 0, 0 },
      '{ 0, 0, 0, 1, 1, 1, 6, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 6, 1, 1, 1, 0, 0, 0 },
      '{ 0, 0, 0, 1, 1, 1, 6, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 6, 1, 1, 1, 0, 0, 0 },
      '{ 0, 0, 0, 1, 1, 6, 6, 1, 1, 1, 1, 1, 6, 1, 6, 1, 1, 1, 1, 1, 6, 6, 1, 1, 0, 0, 0 },
      '{ 0, 0, 1, 1, 1, 6, 1, 6, 6, 6, 6, 6, 1, 1, 1, 6, 6, 6, 6, 6, 1, 6, 1, 1, 1, 0, 0 }, 
      '{ 0, 0, 1, 1, 6, 1, 1, 1, 1, 1, 1, 1, 1, 11, 1, 1, 1, 1, 1, 1, 1, 1, 6, 1, 1, 0, 0 },
      '{ 0, 0, 1, 1, 6, 1, 1, 1, 1, 1, 6, 1, 1, 1, 1, 1, 6, 1, 1, 1, 1, 1, 6, 1, 1, 0, 0 },
      '{ 0, 0, 1, 6, 1, 6, 1, 1, 1, 6, 1, 1, 6, 1, 6, 1, 1, 6, 1, 1, 1, 6, 1, 6, 1, 0, 0 },
      '{ 0, 1, 1, 6, 1, 1, 6, 1, 6, 1, 1, 1, 6, 1, 6, 1, 1, 1, 6, 1, 6, 1, 1, 6, 1, 1, 0 },
      '{ 0, 1, 6, 6, 1, 1, 1, 6, 1, 1, 6, 1, 6, 1, 6, 1, 6, 1, 1, 6, 1, 1, 1, 6, 6, 1, 0 },
      '{ 0, 1, 6, 6, 1, 1, 1, 1, 6, 1, 6, 1, 6, 1, 6, 1, 6, 1, 6, 1, 1, 1, 1, 6, 6, 1, 0 },
      '{ 1, 6, 6, 1, 1, 1, 1, 11, 1, 6, 6, 1, 6, 1, 6, 1, 6, 6, 1, 11, 1, 1, 1, 1, 6, 6, 1 }, 
      '{ 1, 6, 6, 1, 1, 1, 1, 1, 1, 1, 6, 6, 6, 6, 6, 6, 6, 1, 1, 1, 1, 1, 1, 1, 6, 6, 1 }, 
      '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0 }
    };


    //1-Shell (16 x 16)
    Oneshell_font <= '{
      '{0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
      '{0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0 },
      '{0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0 },
      '{0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0 },
      '{0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0 },
      '{0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0 },
      '{0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0 },
      '{1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1 },
      '{1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1 },
      '{1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1 }, 
      '{11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11 },
      '{1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1 }, 
      '{0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0 },  
      '{0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0 }, 
      '{0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0 },
      '{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }
    };


  //2-Shell (33 x 16){
   Twoshell_font <= '{ 
     '{0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
     '{0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0 },
     '{0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0 },
     '{0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0 },
     '{0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0 },
     '{0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0 },
     '{0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0 },
     '{1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1 },
     '{1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1 },
     '{1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1, 0, 1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1 },
     '{11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11, 0, 11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11 },
     '{1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1, 0, 1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1 },
     '{0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0, 0, 0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0 },
     '{0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0, 0, 0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0 }, 
     '{0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0 },
     '{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 } 
    };


   //3-Shell (50 x 16)
   Threeshell_font <= '{
   '{0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },
   '{0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0 },
   '{0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0 },
   '{0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 0, 0 },
   '{0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0 },
   '{0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 0 },
   '{0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0 },
   '{1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1 },
   '{1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1 },
   '{1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1, 0, 1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1, 0, 1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1 },
   '{11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11, 0, 11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11, 0, 11, 11, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 11, 11 },
   '{1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1, 0, 1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1, 0, 1, 11, 11, 11, 1, 2, 2, 2, 2, 2, 2, 1, 11, 11, 11, 1 }, 
   '{0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0, 0, 0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0, 0, 0, 1, 1, 11, 11, 1, 1, 1, 1, 1, 1, 11, 11, 1, 1, 0 },
   '{0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0, 0, 0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0, 0, 0, 0, 0, 1, 11, 11, 11, 11, 11, 11, 11, 11, 1, 0, 0, 0 },
   '{0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 11, 11, 11, 11, 1, 1, 0, 0, 0, 0 },
   '{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }    
   };

	//Police Car (28 x 12)
	policecar_font <= '{
	'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4,10, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,11, 6, 6, 6,11, 6, 6, 6,11, 1, 0, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,11, 6, 6, 6, 6,11, 6, 6, 6, 6,11, 1, 0, 0, 0, 0, 0 },  
	'{0, 0, 0, 0, 0, 0, 0, 1, 1, 1,11, 6, 6, 6, 6, 6,11, 6, 6, 6, 6,11,11, 1, 0, 0, 0, 0 },
	'{0, 0, 0, 1, 1, 1, 1,13,13, 1,11,11,11,11,11,11,11,11,11,11,11,11,11, 1, 1, 1, 0, 0 }, 
	'{0, 5, 1,13,13, 1, 1,13,13, 1,11,11,11,11,11,11,11,11,11,11,11,11, 1, 1,13,13, 1, 0 },
	'{5, 3,13,13, 1, 6, 6, 1,13, 1,13,13,13,13,13,13,13,13,13,13,13, 1, 6, 6, 1,13, 3, 5 }, 
	'{0, 1, 1, 1, 6, 6, 6, 6, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 6, 6, 6, 6, 1, 1, 0 },
	'{0, 0, 0, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0 } 
	};

	
	// Truck (25 x 14)
	truck_font <= '{
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 6, 6, 0, 8, 0, 8, 0, 8, 0, 8, 0, 8, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 6, 6, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 6, 6, 6, 6, 6, 6, 6, 0, 8, 0, 8, 0, 8, 0, 8, 0, 8, 0, 0 }, 
	'{ 0, 0,10,10,10,10,13,10,10,10,10,13,13,10,10,10,10,10,10,10,10,10,10, 0, 0 }, 
	'{ 0, 5, 7,10,10,10,13,10,10,10,10,10,13,10,10,10,10,10,10,10,10,10, 7, 3, 0 },
	'{ 0, 5,10,10,10,10,13,13,10,10,10,10,13,10,10,10,10,10,10,10,10,10,10, 3, 0 },
	'{ 0,10,10, 1, 1, 1, 1,13,13,10,10,10,13,10,10,10,10,10, 1, 1, 1, 1,10,10, 0 },
	'{ 6,10, 1, 1, 1, 1, 1, 1,13,13,13,13,13,10,10,10,10, 1, 1, 1, 1, 1, 1,10, 6 },
	'{ 6,10, 1, 1, 6, 6, 1, 1,10, 6, 6, 6, 6, 6, 6, 6,10, 1, 1, 6, 6, 1, 1,10, 6 }, 
	'{ 0, 0, 1, 1, 6, 6, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 6, 6, 1, 1, 0, 0 }, 
	'{ 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0 }, 
	'{ 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0 } 
	};


   // Skull (23 x 18)
	skull_font <= '{
	'{0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0 }, 
	'{1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1 }, 
	'{1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1 }, 
	'{0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0 },
	'{0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0 },  
	'{0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }, 
	'{0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }, 
	'{0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0 },
	'{0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0 }, 
	'{1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1 }, 
	'{1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1 }, 
	'{0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0 } 
	};
	
	
	
	
	end
endmodule

