module digitfont( input logic Clk,
               	    // from right to left
               	    input logic digit,  	
					output logic [0:13][0:13][0:5] font 
				  );


logic [0:13][0:13][0:5] zero_font ;  
logic [0:13][0:13][0:5] one_font ; 
logic [0:13][0:13][0:5] two_font ; 
logic [0:13][0:13][0:5] three_font ;  
logic [0:13][0:13][0:5] four_font ;  
logic [0:13][0:13][0:5] five_font ; 
logic [0:13][0:13][0:5] six_font ;
logic [0:13][0:13][0:5] seven_font ; 
logic [0:13][0:13][0:5] eight_font ; 
logic [0:13][0:13][0:5] nine_font ; 



// assign the font values
always_comb
begin
	zero_font <= '{
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{0, 0, 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	'{0, 0, 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	'{0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }
	};

	one_font<='{
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }
	};

	two_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }
	};

	three_font<='{
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	four_font<='{
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	};


	five_font<='{
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	 '{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	};


	six_font<='{
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	seven_font<='{
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 },
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }, 
	'{ 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0 }
	};

	eight_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2 },  
	'{ 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2 },   
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }, 
	'{ 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2 },
	'{ 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 }
	};

	nine_font<='{
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },  
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2 }, 
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 },
	'{ 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0 }, 
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 },
	'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0 }
	};
end 

//output the value

always_comb
begin
	case (digit)
		0 : 
			begin 	
				font = zero_font ; 
			end	
		
		1 : 
			begin 	
				font = one_font ; 
			end	

		2 : 
			begin 	
				font = two_font ; 
			end	

		3 : 
			begin 	
				font = three_font ; 
			end		

		4 : 
			begin 	
				font = four_font ; 
			end		

		5 : 
			begin 	
				font = five_font ; 
			end	

		6 : 
			begin 	
				font = six_font ; 
			end

		7 : 
			begin 	
				font = seven_font ; 
			end		

		8 : 
			begin 	
				font = eight_font ; 
			end	
		
		9 : 
			begin 	
				font = nine_font ; 
			end	

		default : 
			begin      
				font = zero_font ; 
			end 	
		
	endcase	



end

endmodule





endmodule 
